----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:52:12 04/05/2020 
-- Design Name: 
-- Module Name:    ROM_IR - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ROM_IR is
	port(
		address : in std_logic_vector(7 downto 0);
		instruction : out std_logic_vector(7 downto 0);
		data : out std_logic_vector(7 downto 0));
end ROM_IR;

architecture Behavioral of ROM_IR is

type ROM  is array (0 to 255) of std_logic_vector(7 downto 0);

constant ROM_TABLE : ROM := 
      ("00000001","00001010","00001001","00000000", -- 0 
		 "00000001","00001000","00001000","00000010", -- 4
		 "00001100","00111000","00000001","00011100", -- 8
		 "00001000","01100100","00000000","00000000", -- 12
		 "00000000","00000000","00000000","00000000", -- 16
		 "00000000","00000000","00000000","00000000", -- 20
		 "00000000","00000000","00000000","00000000", -- 24
		 "00000000","00000000","00000000","00000000", -- 28
		 "00000000","00000000","00000000","00000000", -- 32
		 "00000000","00000000","00000000","00000000", -- 36
		 "00000000","00000000","00000000","00000000", -- 40
		 "00000000","00000000","00000000","00000000", -- 44
		 "00000000","00000000","00000000","00000000", -- 48
		 "00000000","00000000","00000000","00000000", -- 52
		 "00000001","00011100","00000111","01100001", -- 56
		 "00000000","00000000","00000000","00000000", -- 60
		 "00000000","00000000","00000000","00000000", -- 64 
		 "00000000","00000000","00000000","00000000", -- 68
		 "00000000","00000000","00000000","00000000", -- 72
		 "00000000","00000000","00000000","00000000", -- 76
		 "00000000","00000000","00000000","00000000", -- 80
		 "00000000","00000000","00000000","00000000", -- 84
		 "00000000","00000000","00000000","00000000", -- 88
		 "00000000","00000000","00000000","00000000", -- 92
		 "00000000","00000000","00000000","00000000", -- 96 
		 "00000000","00000000","00000000","00000000", -- 100
		 "00000000","00000000","00000000","00000000", -- 104
		 "00000000","00000000","00000000","00000000", -- 108
		 "00000000","00000000","00000000","00000000", -- 112
		 "00000000","00000000","00000000","00000000", -- 116
		 "00000000","00000000","00000000","00000000", -- 120
		 "00000000","00000000","00000000","00000000", -- 124
		 "00000000","00000000","00000000","00000000", -- 128
		 "00000000","00000000","00000000","00000000", -- 132
		 "00000000","00000000","00000000","00000000", -- 136
		 "00000000","00000000","00000000","00000000", -- 140
		 "00000000","00000000","00000000","00000000", -- 144
		 "00000000","00000000","00000000","00000000", -- 148
		 "00000000","00000000","00000000","00000000", -- 152
		 "00000000","00000000","00000000","00000000", -- 156
		 "00000000","00000000","00000000","00000000", -- 160
		 "00000000","00000000","00000000","00000000", -- 164
		 "00000000","00000000","00000000","00000000", -- 168
		 "00000000","00000000","00000000","00000000", -- 172
		 "00000000","00000000","00000000","00000000", -- 176
		 "00000000","00000000","00000000","00000000", -- 180
		 "00000000","00000000","00000000","00000000", -- 184
		 "00000000","00000000","00000000","00000000", -- 188
		 "00000000","00000000","00000000","00000000", -- 192
		 "00000000","00000000","00000000","00000000", -- 196
		 "00000000","00000000","00000000","00000000", -- 200
		 "00000000","00000000","00000000","00000000", -- 204
		 "00000000","00000000","00000000","00000000", -- 208
		 "00000000","00000000","00000000","00000000", -- 212
		 "00000000","00000000","00000000","00000000", -- 216
		 "00000000","00000000","00000000","00000000", -- 220
		 "00000000","00000000","00000000","00000000", -- 224
		 "00000000","00000000","00000000","00000000", -- 228
		 "00000000","00000000","00000000","00000000", -- 232
		 "00000000","00000000","00000000","00000000", -- 236
		 "00000000","00000000","00000000","00000000", -- 240
		 "00000000","00000000","00000000","00000000", -- 244
		 "00000000","00000000","00000000","00000000", -- 248
		 "00000000","00000000","00000000","00000000");-- 252
		 	 
begin

	process(address)
	
		variable ROMValue1 : std_logic_vector(7 downto 0);
		variable ROMValue2 : std_logic_vector(7 downto 0);
		
			begin
		
				ROMValue1 := ROM_TABLE(conv_integer(address));  -- read ROM 
				ROMValue2 := ROM_TABLE(conv_integer((address)+1));  -- read ROM 
				
				instruction <= ROMValue1;
				data <= ROMValue2;
		
		end process;
	


end Behavioral;

